`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/17/2022 01:40:27 PM
// Design Name: 
// Module Name: clk_div_2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module clk_div_2(
    input clk,
    output slow_clk
    );
    
    //  creates a 50% duty cycle clock.
    //  period 2s, so 1s on, 1s off
    
endmodule
